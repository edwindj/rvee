module r

pub struct IntegerVector {
	sexp C.SEXP
}
